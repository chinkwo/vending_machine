// ************************Declaration***************************************
// File name: key_ctrl.v
// Author: YuZhengguo
// Date: 2017/6/15 8:39:57
// Version Number: 1.0
// Abstract:
// Modification history:(including time, version, author and abstract)
// 2017-06-01 00:00 version 1.0 xxx
// Abstract: Initial
// *********************************end**************************************
module key_ctrl  (
							sclk,              // ������������ʱ��: 50Mhz
							rst_n,            // �����������븴λ����
							key_in,           // ���밴���ź�(KEY1~KEY4)
							flag_key				//	��������ź�(KEY1~KEY4)
						);

//===========================================================================
// PORT declarations
//===========================================================================						
input        sclk; 
input        rst_n;
input  [3:0] key_in;
output [3:0] flag_key;

//�Ĵ�������
reg [19:0] count;
reg [3:0] key_scan; //����ɨ��ֵKEY

//===========================================================================
// ��������ֵ��20msɨ��һ��,����Ƶ��С�ڰ���ë��Ƶ�ʣ��൱���˳����˸�Ƶë���źš�
//===========================================================================
always @(posedge sclk or negedge rst_n)     //���ʱ�ӵ������غ͸�λ���½���
begin
   if(!rst_n)                //��λ�źŵ���Ч
      count <= 20'd0;        //��������0
   else
      begin
         if(count ==20'd999_999)   //20msɨ��һ�ΰ���,20ms����(50M/50-1=999_999)
            begin
               count <= 20'b0;     //�������Ƶ�20ms������������
               key_scan <= key_in; //�������������ƽ
            end
         else
            count <= count + 20'b1; //��������1
     end
end
//===========================================================================
// �����ź�����һ��ʱ�ӽ���
//===========================================================================
reg [3:0] key_scan_r;
always @(posedge sclk)
    key_scan_r <= key_scan;       
    
wire [3:0] flag_key = key_scan_r[3:0] & (~key_scan[3:0]);  //����⵽�������½��ر仯ʱ������ð��������£�������Ч 
		
endmodule